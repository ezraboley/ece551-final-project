module digital_core_tb();


